LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

package const_logic is
	constant op_mem : std_logic_vector := "000";
	constant op_arith : std_logic_vector := "001";
	constant op_cmp : std_logic_vector := "010";
	constant op_mul : std_logic_vector := "011";
	constant op_sys : std_logic_vector := "111";	
	
	constant f_mem_movi : std_logic_vector := "00000";
	constant f_mem_movhi : std_logic_vector := "00001";
	constant f_mem_jump : std_logic_vector := "00010";
	
	constant f_arith_and : std_logic_vector := "00000";
	constant f_arith_or : std_logic_vector := "00001";
	constant f_arith_xor : std_logic_vector := "00010";
	constant f_arith_not : std_logic_vector := "00011";
	constant f_arith_add : std_logic_vector := "00100";
	constant f_arith_sub : std_logic_vector := "00101";
	constant f_arith_sha : std_logic_vector := "00110";
	constant f_arith_shl : std_logic_vector := "00111";
	
	constant f_cmp_lt : std_logic_vector := "00000";
	constant f_cmp_le : std_logic_vector := "00001";
	constant f_cmp_eq : std_logic_vector := "00011";
	constant f_cmp_ltu : std_logic_vector := "00100";
	constant f_cmp_leu : std_logic_vector := "00101";
	
	constant f_mul_mul : std_logic_vector := "00000";
	constant f_mul_mulh : std_logic_vector := "00001";
	constant f_mul_mulhu : std_logic_vector := "00010";
	constant f_mul_div : std_logic_vector := "00100";
	constant f_mul_divu : std_logic_vector := "00101";
	
	------f de SYSTEM---------------------------------
	constant f_ei : std_logic_vector := "00000";
	constant f_di : std_logic_vector := "00001";
	constant f_reti : std_logic_vector := "00100";
	constant f_rds : std_logic_vector := "01100";
	constant f_wrs : std_logic_vector := "10000";
	constant f_getiid: std_logic_vector := "01000";
	constant f_wrpi : STD_LOGIC_VECTOR := "10100";
	constant f_wrvi : STD_LOGIC_VECTOR := "10101";
	constant f_wrpd : STD_LOGIC_VECTOR := "10110";
	constant f_wrvd : STD_LOGIC_VECTOR := "10111";
	constant f_flush : STD_LOGIC_VECTOR := "11000";
	
	constant invalid : std_logic_vector := x"CACA";
	
end const_logic;